`timescale 1ns/1ns

module quiz6;

integer A, B;

initial begin
	A = -5'sd16 / 4;
	B = 5'd16 / 4;
end

endmodule