module quiz4;

initial begin
	$display("\\S\\\n\nHardware Programming");
end

endmodule