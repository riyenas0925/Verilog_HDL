module ALU (CTRL, NUM, A, B, Y);

input [4:0] NUM;
input [31:0] A, B;
output reg [31:0] Y;

endmodule