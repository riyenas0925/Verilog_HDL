`timescale 1ns/1ns

module quiz1;

wire [3:0] a, b, c;

assign a = 4'b0zz1;
assign b = 4'b10x0;
assign c = 4'b1100;

endmodule